* SPICE3 file created from nor.ext - technology: scmos

.option scale=0.1u

M1000 out in1 gnd gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1001 temp in2 vdd vdd pfet w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1002 out in1 temp vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 out in2 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd out 0.07fF
C1 in1 out 0.02fF
C2 temp out 0.04fF
C3 vdd in2 0.07fF
C4 vdd in1 0.07fF
C5 vdd temp 0.12fF
C6 in2 in1 0.06fF
C7 out gnd 0.09fF
C8 in1 gnd 0.20fF
C9 in2 gnd 0.14fF
C10 vdd gnd 0.52fF
