magic
tech scmos
timestamp 1598079838
<< nwell >>
rect -13 -6 19 15
<< ntransistor >>
rect -2 -16 0 -12
rect 6 -24 8 -20
<< ptransistor >>
rect -2 0 0 4
rect 6 0 8 4
<< ndiffusion >>
rect -3 -16 -2 -12
rect 0 -16 1 -12
rect 5 -24 6 -20
rect 8 -24 9 -20
<< pdiffusion >>
rect -3 0 -2 4
rect 0 0 1 4
rect 5 0 6 4
rect 8 0 9 4
<< ndcontact >>
rect -7 -16 -3 -12
rect 1 -16 5 -12
rect 1 -24 5 -20
rect 9 -24 13 -20
<< pdcontact >>
rect -7 0 -3 4
rect 1 0 5 4
rect 9 0 13 4
<< psubstratepcontact >>
rect -7 -24 -3 -20
<< nsubstratencontact >>
rect -7 8 -3 12
<< polysilicon >>
rect -2 4 0 6
rect 6 4 8 6
rect -2 -8 0 0
rect -13 -10 0 -8
rect -2 -12 0 -10
rect -2 -18 0 -16
rect 6 -20 8 0
rect 6 -25 8 -24
rect 6 -27 19 -25
<< metal1 >>
rect -13 8 -7 12
rect -3 8 19 12
rect -7 4 -3 8
rect 1 4 5 5
rect 9 -12 13 0
rect 5 -16 19 -12
rect -7 -20 -3 -16
rect 9 -20 13 -16
rect -3 -24 1 -20
<< labels >>
rlabel metal1 3 10 3 10 5 vdd!
rlabel metal1 -1 -22 -1 -22 1 gnd!
rlabel polysilicon -1 -9 -1 -9 1 in2
rlabel polysilicon 7 -9 7 -9 1 in1
rlabel metal1 16 -14 16 -14 7 out
rlabel pdcontact 3 2 3 2 1 temp
<< end >>
