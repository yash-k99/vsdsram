magic
tech scmos
timestamp 1599365263
<< nwell >>
rect -9 -3 15 18
<< pwell >>
rect -9 -24 15 -3
<< ntransistor >>
rect 2 -13 4 -9
<< ptransistor >>
rect 2 3 4 7
<< ndiffusion >>
rect 1 -13 2 -9
rect 4 -13 5 -9
<< pdiffusion >>
rect 1 3 2 7
rect 4 3 5 7
<< ndcontact >>
rect -3 -13 1 -9
rect 5 -13 9 -9
<< pdcontact >>
rect -3 3 1 7
rect 5 3 9 7
<< psubstratepcontact >>
rect -3 -21 1 -17
<< nsubstratencontact >>
rect -3 11 1 15
<< polysilicon >>
rect 2 7 4 9
rect 2 -9 4 3
rect 2 -15 4 -13
<< polycontact >>
rect -2 -6 2 -2
<< metal1 >>
rect -3 7 1 11
rect -9 -6 -2 -3
rect 5 -4 9 3
rect 5 -7 15 -4
rect 5 -9 9 -7
rect -3 -17 1 -13
<< bb >>
rect -9 -24 15 18
<< labels >>
rlabel metal1 12 -5 12 -5 4 out
rlabel metal1 -6 -4 -6 -4 4 in
rlabel metal1 -1 9 -1 9 1 vdd!
rlabel metal1 -1 -15 -1 -15 1 gnd!
<< end >>
