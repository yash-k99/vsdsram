DFF
.include osu018.lib

M1 clkb clk vdd vdd pfet L=0.2u W=0.4u
M2 clkb clk gnd gnd nfet L=0.2u W=0.4u
M3 1 clk D vdd pfet L=0.2u W=0.4u
M4 1 clkb D gnd nfet L=0.2u W=0.4u 
M5 2 1 vdd vdd pfet L=0.2u W=0.4u
M6 2 1 gnd gnd nfet L=0.2u W=0.4u
M7 3 2 vdd vdd pfet L=0.2u W=0.4u
M8 3 2 gnd gnd nfet L=0.2u W=0.4u
M9 1 clkb 3 vdd pfet L=0.2u W=0.4u
M10 1 clk 3 gnd nfet L=0.2u W=0.4u
M11 4 clkb 2 vdd pfet L=0.2u W=0.4u
M12 4 clk 2 gnd nfet L=0.2u W=0.4u
M13 Q 4 vdd vdd pfet L=0.2u W=0.4u
M14 Q 4 gnd gnd nfet L=0.2u W=0.4u
M15 5 Q vdd vdd pfet L=0.2u W=0.4u
M16 5 Q gnd gnd nfet L=0.2u W=0.4u
M17 4 clk 5 vdd pfet L=0.2u W=0.4u
M18 4 clkb 5 gnd nfet L=0.2u W=0.4u

V1 vdd gnd dc 1.8V
V2 D gnd pulse 0 1.8 2.5ns 60ps 60ps 15ns 30ns
V3 clk gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns

.tran 0.1ns 100ns
.control 
run
plot V(Q) V(D)+2 V(clk)+4
.endc
.end

