magic
tech scmos
timestamp 1598104938
<< nwell >>
rect 13 -52 17 -51
<< polysilicon >>
rect -8 12 -6 21
rect 36 19 53 21
rect -8 10 8 12
rect 6 -9 8 10
rect 6 -11 10 -9
rect 6 -44 8 -11
rect -20 -46 8 -44
rect -20 -66 -18 -46
rect 51 -66 53 19
rect -20 -68 -17 -66
rect 25 -68 53 -66
rect -20 -83 -18 -68
rect -20 -85 8 -83
rect 6 -133 8 -85
rect 51 -91 53 -68
rect 48 -93 53 -91
rect 6 -135 18 -133
rect 51 -134 53 -93
<< polycontact >>
rect 18 -136 22 -132
rect 47 -135 51 -131
<< metal1 >>
rect 10 32 14 35
rect -20 8 10 9
rect -20 7 14 8
rect -20 5 36 7
rect -20 2 -17 5
rect 10 3 36 5
rect 32 2 36 3
rect -35 -24 -31 -22
rect -38 -27 -31 -24
rect -38 -89 -34 -27
rect -21 -50 -18 -22
rect -3 -24 1 -22
rect -3 -27 17 -24
rect -3 -33 1 -27
rect 13 -28 17 -27
rect 32 -28 36 -22
rect 45 -28 49 -27
rect 35 -34 36 -28
rect -21 -53 9 -50
rect 31 -51 34 -48
rect 13 -52 17 -51
rect 33 -52 34 -51
rect 5 -55 9 -53
rect 31 -55 34 -52
rect 9 -58 34 -55
rect 9 -79 26 -78
rect 5 -81 26 -79
rect -23 -84 9 -81
rect -23 -89 -20 -84
rect 2 -107 26 -104
rect -38 -122 -34 -113
rect -24 -114 -21 -113
rect -24 -117 -20 -114
rect -23 -122 -20 -117
rect -6 -122 -2 -117
rect -38 -155 -34 -146
rect -24 -149 -21 -146
rect 2 -149 5 -107
rect 46 -134 47 -131
rect -24 -152 5 -149
rect 22 -155 26 -145
rect -38 -158 26 -155
<< m2contact >>
rect -3 -37 1 -33
rect 45 -52 49 -48
rect -6 -93 -2 -89
rect -6 -117 -2 -113
rect 22 -117 26 -113
rect 46 -149 50 -145
<< metal2 >>
rect -31 -37 -3 -33
rect -31 -85 -27 -37
rect 49 -52 58 -48
rect -31 -88 -2 -85
rect -6 -89 -2 -88
rect -2 -117 22 -113
rect 54 -145 58 -52
rect 50 -149 58 -145
use tg  tg_0
timestamp 1598094814
transform 0 1 21 -1 0 22
box -10 -27 14 15
use inv  inv_0
timestamp 1598077130
transform 0 1 -14 -1 0 -7
box -9 -21 15 18
use tg  tg_1
timestamp 1598094814
transform 0 -1 25 1 0 -12
box -10 -27 14 15
use inv  inv_1
timestamp 1598077130
transform 0 -1 28 1 0 -43
box -9 -21 15 18
use tg  tg_2
timestamp 1598094814
transform 0 -1 -2 -1 0 -65
box -10 -27 14 15
use inv  inv_2
timestamp 1598077130
transform 0 1 -17 -1 0 -98
box -9 -21 15 18
use tg  tg_3
timestamp 1598094814
transform 0 1 33 1 0 -94
box -10 -27 14 15
use inv  inv_3
timestamp 1598077130
transform 0 1 -17 -1 0 -131
box -9 -21 15 18
use inv  inv_4
timestamp 1598077130
transform -1 0 37 0 1 -128
box -9 -21 15 18
<< labels >>
rlabel polysilicon 52 -130 52 -130 7 clk
rlabel metal1 12 34 12 34 5 D
rlabel metal1 12 6 12 6 1 1
rlabel metal1 -20 -30 -20 -30 1 2
rlabel polysilicon 15 -134 15 -134 1 clkb
rlabel metal1 -22 -118 -22 -118 1 Q
rlabel metal1 13 -80 13 -80 1 4
rlabel metal1 -9 -151 -9 -151 1 5
rlabel metal1 34 -25 34 -25 1 3
<< end >>
