Write Driver
.include osu018.lib

.subckt nor2ip in1 in2 out vdd gnd
M1 out in1 gnd gnd nfet L=0.2u W=0.4u
M2 out in2 gnd gnd nfet L=0.2u W=0.4u
M3 out in1 temp vdd pfet L=0.2u W=0.4u
M4 temp in2 vdd vdd pfet L=0.2u W=0.4u
.ends nor2ip

.subckt inv ip op vdd gnd
M1 op ip vdd vdd pfet L=0.2u W=0.4u
M2 op ip gnd gnd nfet L=0.2u W=0.4u
.ends inv

.subckt driver bl blb wb din vdd gnd
xinv1 din dinb vdd gnd inv
xinv2 dinb dinbb vdd gnd inv
xnor2ip1 wb dinb out1 vdd gnd nor2ip
xnor2ip2 wb dinbb out2 vdd gnd nor2ip
M1 blb out1 gnd gnd nfet L=0.2u W=0.4u
M2 bl out2 gnd gnd nfet L=0.2u W=0.4u
.ends driver

M1 bl gnd vdd vdd pfet L=0.2u W=0.2u
M2 blb gnd vdd vdd pfet L=0.2u W=0.2u

V1 vdd gnd dc 1.8V
V2 wb gnd pulse 0 1.8 0 60ps 60ps 2ns 4ns
V3 din gnd pulse 0 1.8 0 60ps 60ps 0.5ns 1ns
xdriver bl blb wb din vdd gnd driver

.tran 0.1p 10n
.control
run
plot V(wb)+6 V(din)+4 V(bl)+2 V(blb)
.endc
.end 
