Sense Amplifier
.include NMOS-180nm.lib
.include PMOS-180nm.lib

.subckt inv ip op vdd gnd
M1 op ip vdd vdd CMOSP L=0.18u W=0.18u
M2 op ip gnd gnd CMOSN L=0.18u W=0.18u
.ends inv

M1 out bl 3 3 CMOSN L=0.18u W=0.18u
M2 2 blb 3 3 CMOSN L=0.18u W=0.18u
M3 out 2 1 1 CMOSP L=0.18u W=0.36u
M4 2 2 1 1 CMOSP L=0.18u W=0.18u
M5 3 rd_en 0 0 CMOSN L=0.18u W=0.36u
xinv out dout 1 0 inv 

Vdd 1 0 dc 1.8v
V2 blb 0 pulse 1.8 0 0 60ps 60ps 1ns 2ns
V3 bl 0 pulse 0 1.8 0 60ps 60ps 1ns 2ns
V4 rd_en 0 pulse 0 1.8 0 60ps 60ps 5ns 10ns

.tran 0.1p 20n
.control
run
plot V(rd_en)
plot V(bl) V(blb)
plot V(dout) 
.endc
.end
