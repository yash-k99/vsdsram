6T SRAM Cell

.include NMOS-180nm.lib
.include PMOS-180nm.lib

*Access Transistors
M1 bl wl q gnd CMOSN L=0.18u W=0.36u
M2 blb wl qb gnd CMOSN L=0.18u W=0.36u
*Inverter 1
M3 q qb vdd vdd CMOSP L=0.18u W=0.36u
M4 q qb gnd gnd CMOSN L=0.18u W=0.72u
*Inverter 2 
M5 qb q vdd vdd CMOSP L=0.18u W=0.36u
M6 qb q gnd gnd CMOSN L=0.18u W=0.72u

V1 vdd gnd dc 1.8v
Vwl wl gnd pulse 0 1.8 0 60ps 60ps 20ns 40ns

*Write Operation
Vbl bl gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns
Vblb blb gnd pulse 1.8 0 0 60ps 60ps 5ns 10ns

.tran 0.1n 100n 
.control
run
plot V(wl)
plot V(bl) V(blb)
plot V(q) V(qb)
.endc
.end
