N-curve

.include osu018.lib

M1 bl wl Q gnd nfet L=0.2u W=0.4u
M2 blb wl Qb gnd nfet L=0.2u W=0.4u
M3 Q Qb gnd gnd nfet L=0.2u W=0.8u
M4 Qb Q gnd gnd nfet L=0.2u W=0.8u
M5 Q Qb vdd vdd pfet L=0.2u W=0.4u
M6 Qb Q vdd vdd pfet L=0.2u W=0.4u

V1 vdd gnd dc 1.8V
Vin Q gnd dc 1.8V
Vwl wl gnd dc 1.8v
Vbl bl gnd dc 1.8v
Vblb blb gnd dc 1.8v

.dc Vin 0 1.8 0.01
.control
run
plot -I(Vin)
.endc
.end
