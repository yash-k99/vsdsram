* SPICE3 file created from cell6T.ext - technology: scmos
.include osu018.lib
.option scale=0.1u

M1000 q qb vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 qb q vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1002 q qb gnd gnd nfet w=8 l=2
+  ad=60 pd=44 as=80 ps=52
M1003 bl wl q gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 qb q gnd gnd nfet w=8 l=2
+  ad=60 pd=44 as=0 ps=0
M1005 blb wl qb gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 qb q 0.26fF
C1 wl bl 0.02fF
C2 qb vdd 0.16fF
C3 qb blb 0.10fF
C4 q vdd 0.22fF
C5 qb bl 0.04fF
C6 q bl 0.04fF
C7 blb gnd 0.02fF
C8 bl gnd 0.03fF
C9 wl gnd 0.21fF
C10 q gnd 0.73fF
C11 qb gnd 0.57fF
C12 vdd gnd 0.64fF

V1 vdd gnd dc 1.8v
Vwl wl gnd pulse 0 1.8 0 60ps 60ps 20ns 40ns
Vbl bl gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns
Vblb blb gnd pulse 1.8 0 0 60ps 60ps 5ns 10ns
.tran 0.1n 100n 
.control
run
plot V(wl)
plot V(bl) V(blb)
plot V(q) V(qb)
.endc
.end
