magic
tech scmos
timestamp 1598094814
<< nwell >>
rect -10 -6 14 15
<< ntransistor >>
rect 1 -16 3 -12
<< ptransistor >>
rect 1 0 3 4
<< ndiffusion >>
rect 0 -16 1 -12
rect 3 -16 4 -12
<< pdiffusion >>
rect 0 0 1 4
rect 3 0 4 4
<< ndcontact >>
rect -4 -16 0 -12
rect 4 -16 8 -12
<< pdcontact >>
rect -4 0 0 4
rect 4 0 8 4
<< psubstratepcontact >>
rect -4 -24 0 -20
<< nsubstratencontact >>
rect -4 8 0 12
<< polysilicon >>
rect 1 4 3 15
rect 1 -2 3 0
rect 1 -12 3 -10
rect 1 -27 3 -16
<< metal1 >>
rect -4 4 0 8
rect -4 -7 0 0
rect -10 -11 0 -7
rect -4 -12 0 -11
rect 4 -7 8 0
rect 4 -11 14 -7
rect 4 -12 8 -11
rect -4 -20 0 -16
<< labels >>
rlabel polysilicon 2 -21 2 -21 1 ncontrol
rlabel polysilicon 2 9 2 9 1 pcontrol
rlabel metal1 -2 -9 -2 -9 1 in
rlabel metal1 10 -9 10 -9 7 out
<< end >>
