* SPICE3 file created from inv.ext - technology: scmos

.option scale=0.1u

M1000 out in gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 out in vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
C0 in out 0.05fF
C1 in vdd 0.13fF
C2 vdd out 0.11fF
C3 out gnd 0.04fF
C4 in gnd 0.11fF
C5 vdd gnd 0.39fF
