magic
tech scmos
timestamp 1598194949
<< polysilicon >>
rect 23 -2 25 0
rect 103 -87 105 -85
<< metal1 >>
rect -10 38 0 41
rect 40 39 50 42
rect 117 38 123 42
rect 43 20 61 24
rect 34 0 39 3
rect 43 0 46 20
rect 54 10 61 14
rect 14 -3 18 0
rect 113 -3 117 25
rect 14 -6 117 -3
rect 14 -101 18 -6
rect 22 -39 24 -36
rect 14 -104 73 -101
rect 80 -104 83 -100
rect 14 -105 77 -104
<< m2contact >>
rect 39 0 43 4
rect 73 -104 77 -100
rect 97 -104 101 -100
rect 80 -119 84 -115
<< metal2 >>
rect 39 -115 43 0
rect 77 -104 97 -100
rect 39 -119 80 -115
use cell6T  cell6T_0
timestamp 1598073530
transform 1 0 13 0 1 55
box -13 -55 27 15
use senseamp  senseamp_0
timestamp 1598076063
transform 1 0 77 0 1 50
box -16 -44 40 20
use writedriver  writedriver_0
timestamp 1598105618
transform 1 0 33 0 1 -54
box -9 -81 120 39
<< labels >>
rlabel metal2 41 -94 41 -94 1 blb
rlabel polysilicon 104 -86 104 -86 1 wb
rlabel metal1 57 12 57 12 1 rd_en
rlabel metal1 120 40 120 40 1 dout
rlabel polysilicon 24 -1 24 -1 1 wl
rlabel metal1 23 -38 23 -38 1 din
rlabel metal1 16 -97 16 -97 1 bl
rlabel metal1 -7 39 -7 39 3 q
rlabel metal1 46 40 46 40 1 qb
<< end >>
