* SPICE3 file created from dff.ext - technology: scmos

.option scale=0.1u

M1000 2 1 vdd vdd pfet w=4 l=2
+  ad=52 pd=42 as=100 ps=90
M1001 5 Q gnd gnd nfet w=4 l=2
+  ad=36 pd=26 as=100 ps=90
M1002 clkb clk vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 4 clkb 5 gnd nfet w=4 l=2
+  ad=64 pd=48 as=0 ps=0
M1004 3 2 gnd gnd nfet w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1005 1 clk 3 gnd nfet w=4 l=2
+  ad=64 pd=48 as=0 ps=0
M1006 4 clk 2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=52 ps=42
M1007 4 clkb 2 vdd pfet w=4 l=2
+  ad=64 pd=48 as=0 ps=0
M1008 1 clkb D gnd nfet w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1009 5 Q vdd vdd pfet w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1010 clkb clk gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 1 clk D vdd pfet w=4 l=2
+  ad=64 pd=48 as=32 ps=24
M1012 Q 4 gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1013 3 2 vdd vdd pfet w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1014 4 clk 5 vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 2 1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 1 clkb 3 vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 Q 4 vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 clkb 3 0.10fF
C1 vdd clk 0.49fF
C2 clkb 5 0.10fF
C3 2 clk 0.01fF
C4 vdd 1 0.22fF
C5 4 5 0.01fF
C6 2 1 0.26fF
C7 vdd clkb 0.34fF
C8 Q 5 0.02fF
C9 clk 1 0.01fF
C10 2 clkb 0.15fF
C11 vdd 4 0.22fF
C12 clk clkb 0.09fF
C13 vdd Q 0.23fF
C14 clk 4 0.01fF
C15 1 clkb 0.56fF
C16 vdd D 0.03fF
C17 clk Q 0.01fF
C18 vdd 3 0.07fF
C19 clkb 4 0.50fF
C20 2 3 0.06fF
C21 vdd 5 0.07fF
C22 clkb Q 0.06fF
C23 1 3 0.01fF
C24 clkb D 0.32fF
C25 4 Q 0.05fF
C26 vdd 2 0.58fF
C27 5 gnd 0.07fF
C28 3 gnd 0.04fF
C29 D gnd 0.03fF
C30 Q gnd 0.23fF
C31 4 gnd 0.39fF
C32 clkb gnd 0.15fF
C33 1 gnd 0.18fF
C34 clk gnd 0.57fF
C35 2 gnd 0.16fF
C36 vdd gnd 3.06fF
