magic
tech scmos
timestamp 1598188025
<< nwell >>
rect -19 -6 145 17
<< ntransistor >>
rect -8 -16 -6 -12
rect 11 -16 13 -12
rect 30 -16 32 -12
rect 46 -16 48 -12
rect 57 -16 59 -12
rect 79 -16 81 -12
rect 98 -16 100 -12
rect 114 -16 116 -12
rect 125 -16 127 -12
<< ptransistor >>
rect -8 0 -6 4
rect 11 0 13 4
rect 30 0 32 4
rect 46 0 48 4
rect 57 0 59 4
rect 79 0 81 4
rect 98 0 100 4
rect 114 0 116 4
rect 125 0 127 4
<< ndiffusion >>
rect -9 -16 -8 -12
rect -6 -16 -5 -12
rect 7 -16 11 -12
rect 13 -16 17 -12
rect 29 -16 30 -12
rect 32 -16 33 -12
rect 45 -16 46 -12
rect 48 -16 49 -12
rect 53 -16 57 -12
rect 59 -16 63 -12
rect 75 -16 79 -12
rect 81 -16 85 -12
rect 97 -16 98 -12
rect 100 -16 101 -12
rect 113 -16 114 -12
rect 116 -16 117 -12
rect 121 -16 125 -12
rect 127 -16 131 -12
<< pdiffusion >>
rect -9 0 -8 4
rect -6 0 -5 4
rect 7 0 11 4
rect 13 0 17 4
rect 29 0 30 4
rect 32 0 33 4
rect 45 0 46 4
rect 48 0 49 4
rect 53 0 57 4
rect 59 0 63 4
rect 75 0 79 4
rect 81 0 85 4
rect 97 0 98 4
rect 100 0 101 4
rect 113 0 114 4
rect 116 0 117 4
rect 121 0 125 4
rect 127 0 131 4
<< ndcontact >>
rect -13 -16 -9 -12
rect -5 -16 -1 -12
rect 3 -16 7 -12
rect 17 -16 21 -12
rect 25 -16 29 -12
rect 33 -16 37 -12
rect 41 -16 45 -12
rect 49 -16 53 -12
rect 63 -16 67 -12
rect 71 -16 75 -12
rect 85 -16 89 -12
rect 93 -16 97 -12
rect 101 -16 105 -12
rect 109 -16 113 -12
rect 117 -16 121 -12
rect 131 -16 135 -12
<< pdcontact >>
rect -13 0 -9 4
rect -5 0 -1 4
rect 3 0 7 4
rect 17 0 21 4
rect 25 0 29 4
rect 33 0 37 4
rect 41 0 45 4
rect 49 0 53 4
rect 63 0 67 4
rect 71 0 75 4
rect 85 0 89 4
rect 93 0 97 4
rect 101 0 105 4
rect 109 0 113 4
rect 117 0 121 4
rect 131 0 135 4
<< psubstratepcontact >>
rect -13 -24 -9 -20
rect 25 -24 29 -20
rect 41 -24 45 -20
rect 93 -24 97 -20
rect 109 -24 113 -20
<< nsubstratencontact >>
rect -13 9 -9 13
rect 25 9 29 13
rect 41 9 45 13
rect 93 9 97 13
rect 109 9 113 13
<< polysilicon >>
rect 46 8 49 12
rect -8 5 13 7
rect -8 4 -6 5
rect 11 4 13 5
rect 30 4 32 6
rect 46 4 48 8
rect 125 6 139 8
rect 57 4 59 6
rect 79 4 81 6
rect 98 4 100 6
rect 114 4 116 6
rect 125 4 127 6
rect -8 -7 -6 0
rect 11 -2 13 0
rect -11 -9 -6 -7
rect -8 -12 -6 -9
rect 30 -5 32 0
rect 26 -7 32 -5
rect 11 -12 13 -11
rect 30 -12 32 -7
rect 46 -5 48 0
rect 57 -1 59 0
rect 79 -1 81 0
rect 42 -7 48 -5
rect 46 -12 48 -7
rect 98 -5 100 0
rect 94 -7 100 -5
rect 57 -12 59 -10
rect 79 -12 81 -10
rect 98 -12 100 -7
rect 114 -5 116 0
rect 125 -2 127 0
rect 110 -7 116 -5
rect 114 -12 116 -7
rect 125 -12 127 -11
rect -8 -25 -6 -16
rect 11 -18 13 -16
rect 30 -18 32 -16
rect 46 -18 48 -16
rect 57 -25 59 -16
rect 79 -25 81 -16
rect 98 -18 100 -16
rect 114 -18 116 -16
rect 125 -18 127 -16
rect 137 -25 139 6
rect -8 -27 139 -25
<< polycontact >>
rect 49 8 54 12
rect -15 -9 -11 -5
rect 10 -11 14 -6
rect 22 -8 26 -4
rect 38 -8 42 -4
rect 56 -6 60 -1
rect 78 -6 82 -1
rect 90 -8 94 -4
rect 106 -8 110 -4
rect 124 -11 128 -6
<< metal1 >>
rect -13 15 113 18
rect -13 13 -9 15
rect -13 4 -9 9
rect 25 13 29 15
rect 25 4 29 9
rect 41 13 45 15
rect 93 13 97 15
rect 41 4 45 9
rect 71 4 75 12
rect 93 4 97 9
rect 109 13 113 15
rect 109 4 113 9
rect -5 -5 -1 0
rect -19 -9 -15 -6
rect -5 -12 -1 -9
rect 3 -12 7 0
rect 17 -4 21 0
rect 33 -4 37 0
rect 17 -8 22 -4
rect 33 -8 38 -4
rect 17 -12 21 -8
rect 33 -12 37 -8
rect 49 -12 53 0
rect -13 -20 -9 -16
rect 63 -12 67 0
rect 71 -12 75 0
rect 85 -4 89 0
rect 101 -4 105 0
rect 85 -8 90 -4
rect 101 -8 106 -4
rect 85 -12 89 -8
rect 101 -12 105 -8
rect 117 -12 121 0
rect 25 -20 29 -16
rect -13 -28 -9 -24
rect 25 -28 29 -24
rect 41 -20 45 -16
rect 131 -12 135 0
rect 93 -20 97 -16
rect 41 -28 45 -24
rect 93 -28 97 -24
rect 109 -20 113 -16
rect 109 -28 113 -24
rect -13 -31 113 -28
<< m2contact >>
rect 67 8 71 12
rect -5 -9 0 -5
rect 17 -20 21 -16
rect 63 -20 67 -16
rect 85 -20 89 -16
rect 131 -20 135 -16
<< metal2 >>
rect 46 8 67 12
rect 56 -5 60 -2
rect 0 -9 128 -5
rect 10 -11 14 -9
rect 124 -11 128 -9
rect 21 -20 63 -16
rect 89 -20 131 -16
<< labels >>
rlabel metal1 -17 -8 -17 -8 3 clk
rlabel metal1 -3 -11 -3 -11 1 clkb
rlabel metal1 5 -10 5 -10 1 D
rlabel metal1 19 -10 19 -10 1 1
rlabel metal1 35 -10 35 -10 1 2
rlabel metal1 51 -10 51 -10 1 3
rlabel metal1 87 -10 87 -10 1 4
rlabel metal1 103 -10 103 -10 1 Q
rlabel metal1 119 -10 119 -10 1 5
rlabel metal1 51 -30 51 -30 1 gnd!
rlabel metal1 43 17 43 17 5 vdd!
<< end >>
