* SPICE3 file created from cell6T.ext - technology: scmos

.option scale=0.1u

M1000 q qb vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 qb q vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1002 q qb gnd gnd nfet w=8 l=2
+  ad=60 pd=44 as=80 ps=52
M1003 bl wl q gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 qb q gnd gnd nfet w=8 l=2
+  ad=60 pd=44 as=0 ps=0
M1005 blb wl qb gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
