* SPICE3 file created from 1bitsram.ext - technology: scmos
.include osu018.lib
.option scale=0.1u

M1000 writedriver_0/inv_1/in din gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 writedriver_0/inv_1/in din vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 writedriver_0/inv_1/out writedriver_0/inv_1/in gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 writedriver_0/inv_1/out writedriver_0/inv_1/in vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 writedriver_0/nor_0/out wb gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 writedriver_0/nor_0/temp writedriver_0/inv_1/in vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 writedriver_0/nor_0/out wb writedriver_0/nor_0/temp vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 writedriver_0/nor_0/out writedriver_0/inv_1/in gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 writedriver_0/nor_1/out writedriver_0/inv_1/out gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 writedriver_0/nor_1/temp wb vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 writedriver_0/nor_1/out writedriver_0/inv_1/out writedriver_0/nor_1/temp vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 writedriver_0/nor_1/out wb gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 bl gnd vdd vdd pfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 blb gnd vdd vdd pfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 bl writedriver_0/nor_1/out gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 blb writedriver_0/nor_0/out gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 q qb vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 qb q vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 q qb gnd gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 bl wl q gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 qb q gnd gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 blb wl qb gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 dout senseamp_0/out vdd vdd pfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 senseamp_0/2 senseamp_0/2 vdd vdd pfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 senseamp_0/out bl senseamp_0/3 gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 senseamp_0/out senseamp_0/2 vdd vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 senseamp_0/2 blb senseamp_0/3 gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 senseamp_0/3 rd_en gnd gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 dout senseamp_0/out gnd gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
C0 wb writedriver_0/inv_1/out 0.07fF
C1 blb writedriver_0/nor_0/out 0.05fF
C2 vdd writedriver_0/nor_1/temp 0.12fF
C3 writedriver_0/inv_1/in writedriver_0/inv_1/out 0.05fF
C4 vdd q 0.22fF
C5 senseamp_0/2 bl 0.01fF
C6 vdd writedriver_0/nor_1/out 0.07fF
C7 vdd senseamp_0/out 0.17fF
C8 bl wl 0.05fF
C9 bl qb 0.09fF
C10 wb writedriver_0/nor_1/out 0.01fF
C11 senseamp_0/3 senseamp_0/out 0.04fF
C12 writedriver_0/nor_0/temp writedriver_0/nor_0/out 0.04fF
C13 vdd blb 0.26fF
C14 senseamp_0/2 vdd 0.27fF
C15 blb rd_en 0.03fF
C16 writedriver_0/inv_1/out writedriver_0/nor_1/out 0.24fF
C17 blb senseamp_0/3 0.08fF
C18 vdd qb 0.20fF
C19 senseamp_0/2 senseamp_0/3 0.14fF
C20 writedriver_0/nor_1/temp writedriver_0/nor_1/out 0.04fF
C21 vdd writedriver_0/nor_0/temp 0.12fF
C22 din vdd 0.15fF
C23 vdd writedriver_0/nor_0/out 0.07fF
C24 bl dout 0.10fF
C25 bl vdd 0.27fF
C26 din writedriver_0/inv_1/in 0.05fF
C27 bl rd_en 0.02fF
C28 q wl 0.06fF
C29 writedriver_0/nor_0/out wb 0.09fF
C30 qb q 0.26fF
C31 vdd dout 0.07fF
C32 senseamp_0/2 blb 0.01fF
C33 blb wl 0.08fF
C34 blb qb 0.22fF
C35 vdd wb 0.16fF
C36 bl q 0.15fF
C37 vdd writedriver_0/inv_1/in 0.59fF
C38 qb wl 0.02fF
C39 bl writedriver_0/nor_1/out 0.11fF
C40 writedriver_0/inv_1/in wb 0.06fF
C41 vdd writedriver_0/inv_1/out 0.39fF
C42 bl senseamp_0/out 0.01fF
C43 rd_en gnd 0.02fF
C44 bl gnd 0.34fF
C45 blb gnd 0.26fF
C46 wl gnd 0.03fF
C47 qb gnd 0.03fF
C48 writedriver_0/nor_1/out gnd 0.21fF
C49 writedriver_0/inv_1/out gnd 0.02fF
C50 wb gnd 0.11fF
C51 writedriver_0/nor_0/out gnd 0.12fF
C52 writedriver_0/inv_1/in gnd 0.05fF
C53 vdd gnd 0.40fF
C54 din gnd 0.02fF

V1 vdd gnd dc 1.8V
Vwl wl gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns
Vq q gnd pulse 0 1.8 0 60ps 60ps 1ns 2ns
Vrd rd_en gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns
Vwb wb gnd dc 1.8V
Vdin din gnd dc 0V

.tran 0.1p 20n
.control
run
plot V(rd_en)+10 V(dout) V(bl)+4 V(blb)+2 V(q)+8 V(qb)+6
.endc
.end
