* SPICE3 file created from tri.ext - technology: scmos

.option scale=0.1u

M1000 out enb 2 vdd pfet w=7 l=2
+  ad=35 pd=24 as=135 ps=60
M1001 out en 3 gnd nfet w=4 l=2
+  ad=20 pd=18 as=120 ps=60
M1002 2 inb vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=84
M1003 inb in gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=120 ps=68
M1004 inb in vdd vdd pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1005 3 inb gnd gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out 2 0.04fF
C1 out enb 0.02fF
C2 vdd inb 0.11fF
C3 vdd in 0.09fF
C4 vdd 2 0.01fF
C5 en inb 0.01fF
C6 en 3 0.04fF
C7 vdd enb 0.18fF
C8 inb in 0.07fF
C9 out vdd 0.12fF
C10 inb enb 0.01fF
C11 out en 0.02fF
C12 in enb 0.01fF
C13 out 3 0.04fF
C14 2 enb 0.03fF
C15 3 gnd 0.01fF
C16 en gnd 0.16fF
C17 out gnd 0.04fF
C18 enb gnd 0.00fF
C19 in gnd 0.11fF
C20 inb gnd 0.15fF
C21 vdd gnd 1.52fF
