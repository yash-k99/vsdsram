Read SNM Calculation

.include osu018.lib

M1 qb1 q1 gnd gnd nfet L=0.2u W=0.8u
M2 qb1 q1 vdd vdd pfet L=0.2u W=0.4u
M5 qb1 vdd vdd gnd nfet L=0.2u W=0.4u
M3 q2 qb2 gnd gnd nfet L=0.2u W=0.8u
M4 q2 qb2 vdd vdd pfet L=0.2u W=0.4u
M6 q2 vdd vdd gnd nfet L=0.2u W=0.4u
V1 vdd gnd 1.8V
V2 q1 gnd dc 1.8V
V3 qb2 gnd dc 1.8V
.dc V2 0 1.8 0.01 V3 0 1.8 0.01

.control
run
plot V(qb1) vs V(q1) V(qb2) vs V(q2) 
.endc
.END
