* SPICE3 file created from writedriver.ext - technology: scmos
.include osu018.lib

M1000 nor_0/in2 inv_0/in gnd gnd nfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0.4p ps=3.6u
M1001 nor_0/in2 inv_0/in vdd vdd pfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1002 inv_0/in din gnd gnd nfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1003 inv_0/in din vdd vdd pfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1004 nor_0/out wb gnd gnd nfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1005 nor_0/temp nor_0/in2 vdd vdd pfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1006 nor_0/out wb nor_0/temp vdd pfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1007 nor_0/out nor_0/in2 gnd gnd nfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1008 nor_1/out wb gnd gnd nfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1009 nor_1/temp inv_0/in vdd vdd pfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1010 nor_1/out wb nor_1/temp vdd pfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1011 nor_1/out inv_0/in gnd gnd nfet w=0.4u l=0.2u
+  ad=0p pd=0u as=0p ps=0u
M1012 bl nor_0/out gnd gnd nfet w=0.4u l=0.2u
+  ad=0.2p pd=1.8u as=0p ps=0u
M1013 blb nor_1/out gnd gnd nfet w=0.4u l=0.2u
+  ad=0.2p pd=1.8u as=0p ps=0u
C0 vdd nor_1/out 0.03fF
C1 nor_1/out nor_1/temp 0.04fF
C2 vdd nor_1/temp 0.06fF
C3 inv_0/in vdd 0.27fF
C4 vdd nor_0/temp 0.06fF
C5 nor_0/out nor_1/out 0.01fF
C6 vdd din 0.13fF
C7 inv_0/in din 0.05fF
C8 vdd nor_0/out 0.03fF
C9 nor_0/temp nor_0/out 0.04fF
C10 nor_0/in2 wb 0.09fF
C11 wb nor_1/out 0.03fF
C12 vdd nor_0/in2 0.19fF
C13 inv_0/in nor_0/in2 0.05fF
C14 vdd wb 0.13fF
C15 inv_0/in wb 0.06fF
C16 nor_0/out wb 0.02fF
C17 bl gnd 0.01fF
C18 blb gnd 0.01fF
C19 nor_1/out gnd 0.21fF
C20 wb gnd 0.43fF
C21 nor_0/out gnd 0.14fF
C22 inv_0/in gnd 0.21fF
C23 din gnd 0.02fF
C24 nor_0/in2 gnd 0.29fF

*Precharge circuit added for simulation purpose only
M1014 bl gnd vdd vdd pfet L=0.2u W=0.3u
M1015 blb gnd vdd vdd pfet L=0.2u W=0.3u

V1 vdd gnd dc 1.8V
V2 wb gnd pulse 0 1.8 0 60ps 60ps 2ns 4ns
V3 din gnd pulse 0 1.8 0 60ps 60ps 0.5ns 1ns

.tran 0.1p 10n
.control
run
plot V(wb)+6 V(din)+4 V(bl)+2 V(blb)
.endc
.end 
