* SPICE3 file created from senseamp.ext - technology: scmos

.option scale=0.1u

M1000 dout out vdd vdd pfet w=3 l=2
+  ad=19 pd=18 as=88 ps=66
M1001 2 2 vdd vdd pfet w=3 l=2
+  ad=19 pd=18 as=0 ps=0
M1002 out bl 3 gnd nfet w=3 l=2
+  ad=19 pd=18 as=88 ps=66
M1003 out 2 vdd vdd pfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 2 blb 3 gnd nfet w=3 l=2
+  ad=19 pd=18 as=0 ps=0
M1005 3 rd_en gnd gnd nfet w=10 l=2
+  ad=0 pd=0 as=69 ps=48
M1006 dout out gnd gnd nfet w=3 l=2
+  ad=19 pd=18 as=0 ps=0
C0 dout bl 0.10fF
C1 blb 3 0.08fF
C2 blb rd_en 0.03fF
C3 bl rd_en 0.02fF
C4 vdd 2 0.27fF
C5 vdd out 0.17fF
C6 vdd dout 0.07fF
C7 vdd blb 0.03fF
C8 vdd bl 0.03fF
C9 2 blb 0.01fF
C10 2 3 0.14fF
C11 2 bl 0.01fF
C12 out 3 0.04fF
C13 out bl 0.01fF
C14 rd_en gnd 0.72fF
C15 3 gnd 0.12fF
C16 bl gnd 0.31fF
C17 blb gnd 0.24fF
C18 dout gnd 0.05fF
C19 out gnd 0.15fF
C20 2 gnd 0.04fF
C21 vdd gnd 1.15fF
