* SPICE3 file created from cell6T.ext - technology: scmos
.include osu018.lib
.option scale=0.1u

M1000 q qb vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 qb q vdd vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1002 q qb gnd gnd nfet w=8 l=2
+  ad=60 pd=44 as=80 ps=52
M1003 bl wl q gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 qb q gnd gnd nfet w=8 l=2
+  ad=60 pd=44 as=0 ps=0
M1005 blb wl qb gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 q wl 0.06fF
C1 qb bl 0.09fF
C2 wl blb 0.08fF
C3 q bl 0.15fF
C4 wl bl 0.05fF
C5 vdd qb 0.20fF
C6 vdd q 0.22fF
C7 vdd blb 0.04fF
C8 qb q 0.26fF
C9 qb blb 0.22fF
C10 qb wl 0.02fF
C11 vdd bl 0.04fF
C12 blb gnd 0.08fF
C13 bl gnd 0.07fF
C14 wl gnd 0.35fF
C15 q gnd 0.41fF
C16 qb gnd 0.32fF
C17 vdd gnd 0.68fF

V1 vdd gnd dc 1.8v
Vwl wl gnd pulse 0 1.8 0 60ps 60ps 20ns 40ns
Vbl bl gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns
Vblb blb gnd pulse 1.8 0 0 60ps 60ps 5ns 10ns
.tran 0.1n 100n 
.control
run
plot V(wl)+8 V(bl)+6 V(blb)+4 V(q)+2 V(qb)
.endc
.end
