magic
tech scmos
timestamp 1599365516
<< pwell >>
rect -36 52 -6 76
rect -26 47 -14 52
rect -12 25 -1 31
rect -7 20 -1 25
<< ntransistor >>
rect -30 63 -26 65
rect -16 63 -12 65
<< ndiffusion >>
rect -30 65 -26 66
rect -16 65 -12 66
rect -30 62 -26 63
rect -16 62 -12 63
<< ndcontact >>
rect -30 66 -26 70
rect -16 66 -12 70
rect -30 58 -26 62
rect -16 58 -12 62
<< psubstratepcontact >>
rect -23 50 -19 54
<< polysilicon >>
rect -35 63 -30 65
rect -26 63 -24 65
rect -18 63 -16 65
rect -12 63 -6 65
rect -35 51 -33 63
rect -25 33 -14 35
rect -25 24 -23 33
rect -9 33 14 35
<< polycontact >>
rect -6 61 -2 65
rect -36 47 -32 51
rect 33 49 37 53
rect -14 32 -9 36
rect -4 5 0 9
<< metal1 >>
rect -30 70 -26 72
rect -16 70 -12 72
rect -26 58 -16 62
rect -23 54 -19 58
rect -6 49 -2 61
rect -36 10 -33 47
rect -6 45 1 49
rect 33 31 37 49
rect 12 28 37 31
rect 0 5 16 9
rect 14 -22 17 -17
<< m2contact >>
rect -30 72 -26 76
rect -16 72 -12 76
rect -14 32 -9 36
<< metal2 >>
rect -30 76 -26 80
rect -30 71 -26 72
rect -16 76 -12 80
rect -16 71 -12 72
rect -36 32 -14 36
rect -9 32 38 36
use nor  nor_0
timestamp 1599365357
transform -1 0 20 0 1 61
box -13 -30 19 15
use inv  inv_0
timestamp 1599365263
transform 0 1 19 1 0 16
box -9 -24 15 18
use nor  nor_1
timestamp 1599365357
transform -1 0 -17 0 -1 -2
box -13 -30 19 15
use inv  inv_1
timestamp 1599365263
transform 0 1 20 1 0 -8
box -9 -24 15 18
<< labels >>
rlabel m2contact -14 73 -14 73 4 bl
rlabel metal1 -21 59 -21 59 4 gnd
rlabel metal1 15 -20 15 -20 4 din
rlabel metal2 19 34 19 34 1 wb
rlabel m2contact -28 73 -28 73 1 blb
<< end >>
