DFF
.include osu018.lib

.subckt tg out in pcontrol ncontrol
M1 out pcontrol in in pfet L=0.2u W=0.4u
M2 out ncontrol in in nfet L=0.2u W=0.4u
.ends tg

.subckt inv out in vdd gnd
M3 out in vdd vdd pfet L=0.2u W=0.4u
M4 out in gnd gnd nfet L=0.2u W=0.4u
.ends inv

.subckt dff D Q clk vdd gnd
xinv1 clkb clk vdd gnd inv 
xtg1 1 D clk clkb tg
xinv2 2 1 vdd gnd inv
xinv3 3 2 vdd gnd inv
xtg2 1 3 clkb clk tg
xtg3 4 2 clkb clk tg
xinv4 Q 4 vdd gnd inv
xinv5 5 Q vdd gnd inv
xtg4 4 5 clk clkb tg
.ends dff

V1 1 0 1.8V
V2 D 0 pulse 0 1.8 0 60ps 60ps 15ns 30ns
V3 clk 0 pulse 0 1.8 0 60ps 60ps 5ns 10ns
xdff D Q clk 1 0 dff
.tran 0.1ns 100ns
.control 
run
plot V(D) 
plot V(Q) 
plot V(clk)
.endc
.end

